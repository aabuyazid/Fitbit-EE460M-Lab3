module FitbitTracker(CLK,pulse,display);

reg [26:0] second_divider;
reg display_change;

reg [7:0] high_activity_counter;


endmodule
